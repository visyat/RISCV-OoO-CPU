module instructionMemory (
    //inputs
    clk, 
    PC, 
    //outputs
    instr, 
    stop
);
    input clk;
    input [31:0] PC; 

    output reg [31:0] instr; 
    output reg stop;

    reg [7:0] instrMem [0:1023];

    initial begin
        for (i=0; i<1024; i++)
            instrMem[i] = 8'b0;
        $readmemh ("instructions.txt", mem) 
        //assumes instructions in hex format; $readmemb for binary
    end

    always @(posedge clk) begin
        if (PC+4 < 1024) begin
            instr = {instrMem[PC],instrMem[PC+1],instrMem[PC+2],instrMem[PC+3]}
            stop = 0;
        end else begin
            instr = 32'b0;
            stop = 1;
        end
    end
endmodule