`timescale 1ns/1ps

module EX_MEM_Reg (
    input           clk,
    input           rstn
);

    always @(posedge clk or negedge rstn) begin
    end

endmodule